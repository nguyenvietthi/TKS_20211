module test();

parameter SIZE=12;

  reg clk;
  reg GO;
  reg signed [SIZE-1:0] storage [0:783]; 
  
  reg we_database;
  reg [SIZE-1:0] dp_database;
  reg [12:0] address_p_database;
  
  reg [9:0] x;
  
  wire [3:0] RESULT;
  TOP TOP(
   .clk                    (clk),
   .GO                     (GO),
   .RESULT                 (RESULT),
   .we_database            (we_database), 
   .dp_database            (dp_database), 
   .address_p_database     (address_p_database-1'b1),
   .STOP                   (STOP)
  );
initial begin
  clk=0;
  address_p_database=0;
  x=0;
  we_database=1;
  #200 GO=1;
end
always #10 clk=~clk;
always @(posedge clk)
   begin
       if (we_database)
       begin
           if (address_p_database<=783) 
               begin
                       dp_database = storage[address_p_database];
                       address_p_database=address_p_database+1'b1;
               end
           else we_database=0;
       end
       if ((x<=28*28)&&(GO)) x=x+1;
       else GO=0;
   if (STOP==1)
   begin
       $display("RESULT: %d",RESULT);
       $finish;
   end
 end
// Precision: 13
// Image size: 28x28
// Answer: 7

initial
begin
	storage[0] =  12'b100011110000; // [0.55859375]
	storage[1] =  12'b100100010000; // [0.56640625]
	storage[2] =  12'b100100110000; // [0.57421875]
	storage[3] =  12'b100101010000; // [0.58203125]
	storage[4] =  12'b100101110000; // [0.58984375]
	storage[5] =  12'b100110000000; // [0.59375]
	storage[6] =  12'b100110100000; // [0.6015625]
	storage[7] =  12'b100110110000; // [0.60546875]
	storage[8] =  12'b100111010000; // [0.61328125]
	storage[9] =  12'b100111100000; // [0.6171875]
	storage[10] =  12'b101000000000; // [0.625]
	storage[11] =  12'b101000000000; // [0.625]
	storage[12] =  12'b101000010000; // [0.62890625]
	storage[13] =  12'b101000010000; // [0.62890625]
	storage[14] =  12'b101000010000; // [0.62890625]
	storage[15] =  12'b101000000000; // [0.625]
	storage[16] =  12'b101000000000; // [0.625]
	storage[17] =  12'b100111100000; // [0.6171875]
	storage[18] =  12'b100111000000; // [0.609375]
	storage[19] =  12'b100110010000; // [0.59765625]
	storage[20] =  12'b100101010000; // [0.58203125]
	storage[21] =  12'b100011110000; // [0.55859375]
	storage[22] =  12'b100011010000; // [0.55078125]
	storage[23] =  12'b100100110000; // [0.57421875]
	storage[24] =  12'b100101110000; // [0.58984375]
	storage[25] =  12'b100110000000; // [0.59375]
	storage[26] =  12'b100101110000; // [0.58984375]
	storage[27] =  12'b100101010000; // [0.58203125]
	storage[28] =  12'b100100010000; // [0.56640625]
	storage[29] =  12'b100100110000; // [0.57421875]
	storage[30] =  12'b100101010000; // [0.58203125]
	storage[31] =  12'b100101110000; // [0.58984375]
	storage[32] =  12'b100110000000; // [0.59375]
	storage[33] =  12'b100110010000; // [0.59765625]
	storage[34] =  12'b100110010000; // [0.59765625]
	storage[35] =  12'b100110100000; // [0.6015625]
	storage[36] =  12'b100110110000; // [0.60546875]
	storage[37] =  12'b100111000000; // [0.609375]
	storage[38] =  12'b100111010000; // [0.61328125]
	storage[39] =  12'b100111010000; // [0.61328125]
	storage[40] =  12'b100111010000; // [0.61328125]
	storage[41] =  12'b100111000000; // [0.609375]
	storage[42] =  12'b100110100000; // [0.6015625]
	storage[43] =  12'b100101110000; // [0.58984375]
	storage[44] =  12'b100101010000; // [0.58203125]
	storage[45] =  12'b100100010000; // [0.56640625]
	storage[46] =  12'b100010010000; // [0.53515625]
	storage[47] =  12'b100000000000; // [0.5]
	storage[48] =  12'b011101100000; // [0.4609375]
	storage[49] =  12'b011011000000; // [0.421875]
	storage[50] =  12'b011100000000; // [0.4375]
	storage[51] =  12'b100000010000; // [0.50390625]
	storage[52] =  12'b100100110000; // [0.57421875]
	storage[53] =  12'b100110000000; // [0.59375]
	storage[54] =  12'b100101110000; // [0.58984375]
	storage[55] =  12'b100101100000; // [0.5859375]
	storage[56] =  12'b100100100000; // [0.5703125]
	storage[57] =  12'b100101000000; // [0.578125]
	storage[58] =  12'b100101010000; // [0.58203125]
	storage[59] =  12'b100101110000; // [0.58984375]
	storage[60] =  12'b100101110000; // [0.58984375]
	storage[61] =  12'b100100110000; // [0.57421875]
	storage[62] =  12'b100010010000; // [0.53515625]
	storage[63] =  12'b100001100000; // [0.5234375]
	storage[64] =  12'b100010010000; // [0.53515625]
	storage[65] =  12'b100010010000; // [0.53515625]
	storage[66] =  12'b100001110000; // [0.52734375]
	storage[67] =  12'b100001000000; // [0.515625]
	storage[68] =  12'b100000000000; // [0.5]
	storage[69] =  12'b011111000000; // [0.484375]
	storage[70] =  12'b011110000000; // [0.46875]
	storage[71] =  12'b011101010000; // [0.45703125]
	storage[72] =  12'b011011110000; // [0.43359375]
	storage[73] =  12'b011010010000; // [0.41015625]
	storage[74] =  12'b011000100000; // [0.3828125]
	storage[75] =  12'b010110100000; // [0.3515625]
	storage[76] =  12'b010100110000; // [0.32421875]
	storage[77] =  12'b010100010000; // [0.31640625]
	storage[78] =  12'b010110110000; // [0.35546875]
	storage[79] =  12'b011101000000; // [0.453125]
	storage[80] =  12'b100011100000; // [0.5546875]
	storage[81] =  12'b100110000000; // [0.59375]
	storage[82] =  12'b100110010000; // [0.59765625]
	storage[83] =  12'b100101110000; // [0.58984375]
	storage[84] =  12'b100100110000; // [0.57421875]
	storage[85] =  12'b100101000000; // [0.578125]
	storage[86] =  12'b100101100000; // [0.5859375]
	storage[87] =  12'b100101110000; // [0.58984375]
	storage[88] =  12'b100101100000; // [0.5859375]
	storage[89] =  12'b100011000000; // [0.546875]
	storage[90] =  12'b011010100000; // [0.4140625]
	storage[91] =  12'b010111000000; // [0.359375]
	storage[92] =  12'b010110100000; // [0.3515625]
	storage[93] =  12'b010110010000; // [0.34765625]
	storage[94] =  12'b010110010000; // [0.34765625]
	storage[95] =  12'b010110010000; // [0.34765625]
	storage[96] =  12'b010110010000; // [0.34765625]
	storage[97] =  12'b010110010000; // [0.34765625]
	storage[98] =  12'b010110010000; // [0.34765625]
	storage[99] =  12'b010110100000; // [0.3515625]
	storage[100] =  12'b010110010000; // [0.34765625]
	storage[101] =  12'b010110000000; // [0.34375]
	storage[102] =  12'b010101000000; // [0.328125]
	storage[103] =  12'b010011110000; // [0.30859375]
	storage[104] =  12'b010010100000; // [0.2890625]
	storage[105] =  12'b010001100000; // [0.2734375]
	storage[106] =  12'b010101000000; // [0.328125]
	storage[107] =  12'b011100100000; // [0.4453125]
	storage[108] =  12'b100011110000; // [0.55859375]
	storage[109] =  12'b100110100000; // [0.6015625]
	storage[110] =  12'b100110100000; // [0.6015625]
	storage[111] =  12'b100110010000; // [0.59765625]
	storage[112] =  12'b100101010000; // [0.58203125]
	storage[113] =  12'b100101100000; // [0.5859375]
	storage[114] =  12'b100101110000; // [0.58984375]
	storage[115] =  12'b100110000000; // [0.59375]
	storage[116] =  12'b100101100000; // [0.5859375]
	storage[117] =  12'b100011000000; // [0.546875]
	storage[118] =  12'b011010010000; // [0.41015625]
	storage[119] =  12'b010100010000; // [0.31640625]
	storage[120] =  12'b010011010000; // [0.30078125]
	storage[121] =  12'b010011000000; // [0.296875]
	storage[122] =  12'b010011110000; // [0.30859375]
	storage[123] =  12'b010101010000; // [0.33203125]
	storage[124] =  12'b010110100000; // [0.3515625]
	storage[125] =  12'b011000000000; // [0.375]
	storage[126] =  12'b011001100000; // [0.3984375]
	storage[127] =  12'b011010110000; // [0.41796875]
	storage[128] =  12'b011011110000; // [0.43359375]
	storage[129] =  12'b011101000000; // [0.453125]
	storage[130] =  12'b011101000000; // [0.453125]
	storage[131] =  12'b011001100000; // [0.3984375]
	storage[132] =  12'b010011110000; // [0.30859375]
	storage[133] =  12'b010010010000; // [0.28515625]
	storage[134] =  12'b010110110000; // [0.35546875]
	storage[135] =  12'b011110110000; // [0.48046875]
	storage[136] =  12'b100101010000; // [0.58203125]
	storage[137] =  12'b100111000000; // [0.609375]
	storage[138] =  12'b100111000000; // [0.609375]
	storage[139] =  12'b100110110000; // [0.60546875]
	storage[140] =  12'b100101010000; // [0.58203125]
	storage[141] =  12'b100101110000; // [0.58984375]
	storage[142] =  12'b100110000000; // [0.59375]
	storage[143] =  12'b100110010000; // [0.59765625]
	storage[144] =  12'b100110000000; // [0.59375]
	storage[145] =  12'b100100100000; // [0.5703125]
	storage[146] =  12'b011111000000; // [0.484375]
	storage[147] =  12'b011001010000; // [0.39453125]
	storage[148] =  12'b011001000000; // [0.390625]
	storage[149] =  12'b011010100000; // [0.4140625]
	storage[150] =  12'b011101000000; // [0.453125]
	storage[151] =  12'b011111010000; // [0.48828125]
	storage[152] =  12'b100001010000; // [0.51953125]
	storage[153] =  12'b100011010000; // [0.55078125]
	storage[154] =  12'b100100100000; // [0.5703125]
	storage[155] =  12'b100101010000; // [0.58203125]
	storage[156] =  12'b100101110000; // [0.58984375]
	storage[157] =  12'b100101100000; // [0.5859375]
	storage[158] =  12'b100011110000; // [0.55859375]
	storage[159] =  12'b011101000000; // [0.453125]
	storage[160] =  12'b010101000000; // [0.328125]
	storage[161] =  12'b010100010000; // [0.31640625]
	storage[162] =  12'b011010110000; // [0.41796875]
	storage[163] =  12'b100010100000; // [0.5390625]
	storage[164] =  12'b100110110000; // [0.60546875]
	storage[165] =  12'b100111100000; // [0.6171875]
	storage[166] =  12'b100111100000; // [0.6171875]
	storage[167] =  12'b100111000000; // [0.609375]
	storage[168] =  12'b100101000000; // [0.578125]
	storage[169] =  12'b100101110000; // [0.58984375]
	storage[170] =  12'b100110010000; // [0.59765625]
	storage[171] =  12'b100110100000; // [0.6015625]
	storage[172] =  12'b100110110000; // [0.60546875]
	storage[173] =  12'b100110100000; // [0.6015625]
	storage[174] =  12'b100101100000; // [0.5859375]
	storage[175] =  12'b100100100000; // [0.5703125]
	storage[176] =  12'b100101000000; // [0.578125]
	storage[177] =  12'b100110010000; // [0.59765625]
	storage[178] =  12'b100111010000; // [0.61328125]
	storage[179] =  12'b101000000000; // [0.625]
	storage[180] =  12'b101000110000; // [0.63671875]
	storage[181] =  12'b101001010000; // [0.64453125]
	storage[182] =  12'b101001010000; // [0.64453125]
	storage[183] =  12'b101001100000; // [0.6484375]
	storage[184] =  12'b101001010000; // [0.64453125]
	storage[185] =  12'b100111110000; // [0.62109375]
	storage[186] =  12'b100100010000; // [0.56640625]
	storage[187] =  12'b011100100000; // [0.4453125]
	storage[188] =  12'b010101110000; // [0.33984375]
	storage[189] =  12'b010111000000; // [0.359375]
	storage[190] =  12'b011111000000; // [0.484375]
	storage[191] =  12'b100101110000; // [0.58984375]
	storage[192] =  12'b100111110000; // [0.62109375]
	storage[193] =  12'b101000010000; // [0.62890625]
	storage[194] =  12'b101000000000; // [0.625]
	storage[195] =  12'b100111100000; // [0.6171875]
	storage[196] =  12'b100101100000; // [0.5859375]
	storage[197] =  12'b100110000000; // [0.59375]
	storage[198] =  12'b100110100000; // [0.6015625]
	storage[199] =  12'b100110110000; // [0.60546875]
	storage[200] =  12'b100111010000; // [0.61328125]
	storage[201] =  12'b100111100000; // [0.6171875]
	storage[202] =  12'b100111110000; // [0.62109375]
	storage[203] =  12'b101000000000; // [0.625]
	storage[204] =  12'b101000100000; // [0.6328125]
	storage[205] =  12'b101001000000; // [0.640625]
	storage[206] =  12'b101001100000; // [0.6484375]
	storage[207] =  12'b101001110000; // [0.65234375]
	storage[208] =  12'b101010100000; // [0.6640625]
	storage[209] =  12'b101010100000; // [0.6640625]
	storage[210] =  12'b101010100000; // [0.6640625]
	storage[211] =  12'b101010100000; // [0.6640625]
	storage[212] =  12'b101010010000; // [0.66015625]
	storage[213] =  12'b101000000000; // [0.625]
	storage[214] =  12'b100011100000; // [0.5546875]
	storage[215] =  12'b011011010000; // [0.42578125]
	storage[216] =  12'b010110100000; // [0.3515625]
	storage[217] =  12'b011010000000; // [0.40625]
	storage[218] =  12'b100010010000; // [0.53515625]
	storage[219] =  12'b100111010000; // [0.61328125]
	storage[220] =  12'b101000100000; // [0.6328125]
	storage[221] =  12'b101000100000; // [0.6328125]
	storage[222] =  12'b101000010000; // [0.62890625]
	storage[223] =  12'b100111110000; // [0.62109375]
	storage[224] =  12'b100101100000; // [0.5859375]
	storage[225] =  12'b100110000000; // [0.59375]
	storage[226] =  12'b100110100000; // [0.6015625]
	storage[227] =  12'b100111000000; // [0.609375]
	storage[228] =  12'b100111100000; // [0.6171875]
	storage[229] =  12'b101000000000; // [0.625]
	storage[230] =  12'b101000100000; // [0.6328125]
	storage[231] =  12'b101000110000; // [0.63671875]
	storage[232] =  12'b101001010000; // [0.64453125]
	storage[233] =  12'b101001100000; // [0.6484375]
	storage[234] =  12'b101010010000; // [0.66015625]
	storage[235] =  12'b101010100000; // [0.6640625]
	storage[236] =  12'b101010110000; // [0.66796875]
	storage[237] =  12'b101011010000; // [0.67578125]
	storage[238] =  12'b101011000000; // [0.671875]
	storage[239] =  12'b101011000000; // [0.671875]
	storage[240] =  12'b101010010000; // [0.66015625]
	storage[241] =  12'b100111110000; // [0.62109375]
	storage[242] =  12'b100001110000; // [0.52734375]
	storage[243] =  12'b011001110000; // [0.40234375]
	storage[244] =  12'b010111010000; // [0.36328125]
	storage[245] =  12'b011101100000; // [0.4609375]
	storage[246] =  12'b100101000000; // [0.578125]
	storage[247] =  12'b101000000000; // [0.625]
	storage[248] =  12'b101000110000; // [0.63671875]
	storage[249] =  12'b101000100000; // [0.6328125]
	storage[250] =  12'b101000010000; // [0.62890625]
	storage[251] =  12'b100111110000; // [0.62109375]
	storage[252] =  12'b100101100000; // [0.5859375]
	storage[253] =  12'b100110010000; // [0.59765625]
	storage[254] =  12'b100110110000; // [0.60546875]
	storage[255] =  12'b100111010000; // [0.61328125]
	storage[256] =  12'b100111110000; // [0.62109375]
	storage[257] =  12'b101000010000; // [0.62890625]
	storage[258] =  12'b101000110000; // [0.63671875]
	storage[259] =  12'b101001100000; // [0.6484375]
	storage[260] =  12'b101001110000; // [0.65234375]
	storage[261] =  12'b101010000000; // [0.65625]
	storage[262] =  12'b101010100000; // [0.6640625]
	storage[263] =  12'b101011000000; // [0.671875]
	storage[264] =  12'b101011010000; // [0.67578125]
	storage[265] =  12'b101011010000; // [0.67578125]
	storage[266] =  12'b101011000000; // [0.671875]
	storage[267] =  12'b101010110000; // [0.66796875]
	storage[268] =  12'b101001110000; // [0.65234375]
	storage[269] =  12'b100110000000; // [0.59375]
	storage[270] =  12'b011110110000; // [0.48046875]
	storage[271] =  12'b011000110000; // [0.38671875]
	storage[272] =  12'b011001110000; // [0.40234375]
	storage[273] =  12'b100001010000; // [0.51953125]
	storage[274] =  12'b100110110000; // [0.60546875]
	storage[275] =  12'b101000110000; // [0.63671875]
	storage[276] =  12'b101000110000; // [0.63671875]
	storage[277] =  12'b101000100000; // [0.6328125]
	storage[278] =  12'b101000000000; // [0.625]
	storage[279] =  12'b100111110000; // [0.62109375]
	storage[280] =  12'b100110000000; // [0.59375]
	storage[281] =  12'b100110100000; // [0.6015625]
	storage[282] =  12'b100110110000; // [0.60546875]
	storage[283] =  12'b100111100000; // [0.6171875]
	storage[284] =  12'b101000000000; // [0.625]
	storage[285] =  12'b101000100000; // [0.6328125]
	storage[286] =  12'b101001000000; // [0.640625]
	storage[287] =  12'b101001010000; // [0.64453125]
	storage[288] =  12'b101001110000; // [0.65234375]
	storage[289] =  12'b101010010000; // [0.66015625]
	storage[290] =  12'b101010110000; // [0.66796875]
	storage[291] =  12'b101011000000; // [0.671875]
	storage[292] =  12'b101011100000; // [0.6796875]
	storage[293] =  12'b101011010000; // [0.67578125]
	storage[294] =  12'b101011000000; // [0.671875]
	storage[295] =  12'b101010100000; // [0.6640625]
	storage[296] =  12'b101000000000; // [0.625]
	storage[297] =  12'b100011010000; // [0.55078125]
	storage[298] =  12'b011011100000; // [0.4296875]
	storage[299] =  12'b011000100000; // [0.3828125]
	storage[300] =  12'b011101110000; // [0.46484375]
	storage[301] =  12'b100101000000; // [0.578125]
	storage[302] =  12'b101000010000; // [0.62890625]
	storage[303] =  12'b101001000000; // [0.640625]
	storage[304] =  12'b101001000000; // [0.640625]
	storage[305] =  12'b101000110000; // [0.63671875]
	storage[306] =  12'b101000010000; // [0.62890625]
	storage[307] =  12'b100111110000; // [0.62109375]
	storage[308] =  12'b100110000000; // [0.59375]
	storage[309] =  12'b100110010000; // [0.59765625]
	storage[310] =  12'b100110110000; // [0.60546875]
	storage[311] =  12'b100111100000; // [0.6171875]
	storage[312] =  12'b101000000000; // [0.625]
	storage[313] =  12'b101000100000; // [0.6328125]
	storage[314] =  12'b101001000000; // [0.640625]
	storage[315] =  12'b101001110000; // [0.65234375]
	storage[316] =  12'b101010000000; // [0.65625]
	storage[317] =  12'b101010010000; // [0.66015625]
	storage[318] =  12'b101011000000; // [0.671875]
	storage[319] =  12'b101011010000; // [0.67578125]
	storage[320] =  12'b101011100000; // [0.6796875]
	storage[321] =  12'b101011010000; // [0.67578125]
	storage[322] =  12'b101011000000; // [0.671875]
	storage[323] =  12'b101010000000; // [0.65625]
	storage[324] =  12'b100110010000; // [0.59765625]
	storage[325] =  12'b011111010000; // [0.48828125]
	storage[326] =  12'b011001100000; // [0.3984375]
	storage[327] =  12'b011010000000; // [0.40625]
	storage[328] =  12'b100001110000; // [0.52734375]
	storage[329] =  12'b100111010000; // [0.61328125]
	storage[330] =  12'b101000110000; // [0.63671875]
	storage[331] =  12'b101001100000; // [0.6484375]
	storage[332] =  12'b101001100000; // [0.6484375]
	storage[333] =  12'b101000110000; // [0.63671875]
	storage[334] =  12'b101000010000; // [0.62890625]
	storage[335] =  12'b101000000000; // [0.625]
	storage[336] =  12'b100101110000; // [0.58984375]
	storage[337] =  12'b100110010000; // [0.59765625]
	storage[338] =  12'b100110110000; // [0.60546875]
	storage[339] =  12'b100111100000; // [0.6171875]
	storage[340] =  12'b101000100000; // [0.6328125]
	storage[341] =  12'b101001000000; // [0.640625]
	storage[342] =  12'b101001110000; // [0.65234375]
	storage[343] =  12'b101010000000; // [0.65625]
	storage[344] =  12'b101010100000; // [0.6640625]
	storage[345] =  12'b101010110000; // [0.66796875]
	storage[346] =  12'b101011010000; // [0.67578125]
	storage[347] =  12'b101011100000; // [0.6796875]
	storage[348] =  12'b101011100000; // [0.6796875]
	storage[349] =  12'b101011100000; // [0.6796875]
	storage[350] =  12'b101011000000; // [0.671875]
	storage[351] =  12'b101001000000; // [0.640625]
	storage[352] =  12'b100011100000; // [0.5546875]
	storage[353] =  12'b011011110000; // [0.43359375]
	storage[354] =  12'b011000100000; // [0.3828125]
	storage[355] =  12'b011101000000; // [0.453125]
	storage[356] =  12'b100100100000; // [0.5703125]
	storage[357] =  12'b101000100000; // [0.6328125]
	storage[358] =  12'b101001010000; // [0.64453125]
	storage[359] =  12'b101001110000; // [0.65234375]
	storage[360] =  12'b101001110000; // [0.65234375]
	storage[361] =  12'b101001000000; // [0.640625]
	storage[362] =  12'b101000010000; // [0.62890625]
	storage[363] =  12'b101000000000; // [0.625]
	storage[364] =  12'b100110000000; // [0.59375]
	storage[365] =  12'b100110110000; // [0.60546875]
	storage[366] =  12'b100111100000; // [0.6171875]
	storage[367] =  12'b101000000000; // [0.625]
	storage[368] =  12'b101001000000; // [0.640625]
	storage[369] =  12'b101001010000; // [0.64453125]
	storage[370] =  12'b101010000000; // [0.65625]
	storage[371] =  12'b101010100000; // [0.6640625]
	storage[372] =  12'b101010110000; // [0.66796875]
	storage[373] =  12'b101011000000; // [0.671875]
	storage[374] =  12'b101011010000; // [0.67578125]
	storage[375] =  12'b101011100000; // [0.6796875]
	storage[376] =  12'b101011100000; // [0.6796875]
	storage[377] =  12'b101011010000; // [0.67578125]
	storage[378] =  12'b101010100000; // [0.6640625]
	storage[379] =  12'b100111000000; // [0.609375]
	storage[380] =  12'b100000010000; // [0.50390625]
	storage[381] =  12'b011001100000; // [0.3984375]
	storage[382] =  12'b011001000000; // [0.390625]
	storage[383] =  12'b100000000000; // [0.5]
	storage[384] =  12'b100110110000; // [0.60546875]
	storage[385] =  12'b101001000000; // [0.640625]
	storage[386] =  12'b101001110000; // [0.65234375]
	storage[387] =  12'b101001110000; // [0.65234375]
	storage[388] =  12'b101010000000; // [0.65625]
	storage[389] =  12'b101001010000; // [0.64453125]
	storage[390] =  12'b101000010000; // [0.62890625]
	storage[391] =  12'b100111110000; // [0.62109375]
	storage[392] =  12'b100110100000; // [0.6015625]
	storage[393] =  12'b100111000000; // [0.609375]
	storage[394] =  12'b100111100000; // [0.6171875]
	storage[395] =  12'b101000010000; // [0.62890625]
	storage[396] =  12'b101001000000; // [0.640625]
	storage[397] =  12'b101001010000; // [0.64453125]
	storage[398] =  12'b101010000000; // [0.65625]
	storage[399] =  12'b101010100000; // [0.6640625]
	storage[400] =  12'b101010110000; // [0.66796875]
	storage[401] =  12'b101011010000; // [0.67578125]
	storage[402] =  12'b101011100000; // [0.6796875]
	storage[403] =  12'b101011100000; // [0.6796875]
	storage[404] =  12'b101011100000; // [0.6796875]
	storage[405] =  12'b101010100000; // [0.6640625]
	storage[406] =  12'b101001100000; // [0.6484375]
	storage[407] =  12'b100100110000; // [0.57421875]
	storage[408] =  12'b011101000000; // [0.453125]
	storage[409] =  12'b010111110000; // [0.37109375]
	storage[410] =  12'b011010100000; // [0.4140625]
	storage[411] =  12'b100010000000; // [0.53125]
	storage[412] =  12'b100111000000; // [0.609375]
	storage[413] =  12'b101000110000; // [0.63671875]
	storage[414] =  12'b101001100000; // [0.6484375]
	storage[415] =  12'b101001110000; // [0.65234375]
	storage[416] =  12'b101001110000; // [0.65234375]
	storage[417] =  12'b101001000000; // [0.640625]
	storage[418] =  12'b101000100000; // [0.6328125]
	storage[419] =  12'b100111100000; // [0.6171875]
	storage[420] =  12'b100110010000; // [0.59765625]
	storage[421] =  12'b100110110000; // [0.60546875]
	storage[422] =  12'b100111100000; // [0.6171875]
	storage[423] =  12'b101000100000; // [0.6328125]
	storage[424] =  12'b101000110000; // [0.63671875]
	storage[425] =  12'b101001010000; // [0.64453125]
	storage[426] =  12'b101010000000; // [0.65625]
	storage[427] =  12'b101010100000; // [0.6640625]
	storage[428] =  12'b101011000000; // [0.671875]
	storage[429] =  12'b101011010000; // [0.67578125]
	storage[430] =  12'b101011010000; // [0.67578125]
	storage[431] =  12'b101010110000; // [0.66796875]
	storage[432] =  12'b101001110000; // [0.65234375]
	storage[433] =  12'b101000010000; // [0.62890625]
	storage[434] =  12'b100101110000; // [0.58984375]
	storage[435] =  12'b100000010000; // [0.50390625]
	storage[436] =  12'b011000110000; // [0.38671875]
	storage[437] =  12'b010101010000; // [0.33203125]
	storage[438] =  12'b011000000000; // [0.375]
	storage[439] =  12'b011101000000; // [0.453125]
	storage[440] =  12'b100010100000; // [0.5390625]
	storage[441] =  12'b100111010000; // [0.61328125]
	storage[442] =  12'b101001000000; // [0.640625]
	storage[443] =  12'b101001010000; // [0.64453125]
	storage[444] =  12'b101001010000; // [0.64453125]
	storage[445] =  12'b101001000000; // [0.640625]
	storage[446] =  12'b101000010000; // [0.62890625]
	storage[447] =  12'b100111110000; // [0.62109375]
	storage[448] =  12'b100110010000; // [0.59765625]
	storage[449] =  12'b100111000000; // [0.609375]
	storage[450] =  12'b100111110000; // [0.62109375]
	storage[451] =  12'b101000100000; // [0.6328125]
	storage[452] =  12'b101000110000; // [0.63671875]
	storage[453] =  12'b101001000000; // [0.640625]
	storage[454] =  12'b101001110000; // [0.65234375]
	storage[455] =  12'b101010010000; // [0.66015625]
	storage[456] =  12'b101010100000; // [0.6640625]
	storage[457] =  12'b101010110000; // [0.66796875]
	storage[458] =  12'b101010100000; // [0.6640625]
	storage[459] =  12'b100111010000; // [0.61328125]
	storage[460] =  12'b100001110000; // [0.52734375]
	storage[461] =  12'b011101100000; // [0.4609375]
	storage[462] =  12'b011010010000; // [0.41015625]
	storage[463] =  12'b010111000000; // [0.359375]
	storage[464] =  12'b010011010000; // [0.30078125]
	storage[465] =  12'b010010010000; // [0.28515625]
	storage[466] =  12'b010100000000; // [0.3125]
	storage[467] =  12'b011000010000; // [0.37890625]
	storage[468] =  12'b011111110000; // [0.49609375]
	storage[469] =  12'b100110010000; // [0.59765625]
	storage[470] =  12'b101000100000; // [0.6328125]
	storage[471] =  12'b101001000000; // [0.640625]
	storage[472] =  12'b101001000000; // [0.640625]
	storage[473] =  12'b101000100000; // [0.6328125]
	storage[474] =  12'b101000000000; // [0.625]
	storage[475] =  12'b100111100000; // [0.6171875]
	storage[476] =  12'b100110010000; // [0.59765625]
	storage[477] =  12'b100111000000; // [0.609375]
	storage[478] =  12'b100111110000; // [0.62109375]
	storage[479] =  12'b101000010000; // [0.62890625]
	storage[480] =  12'b101000100000; // [0.6328125]
	storage[481] =  12'b101001000000; // [0.640625]
	storage[482] =  12'b101001100000; // [0.6484375]
	storage[483] =  12'b101001110000; // [0.65234375]
	storage[484] =  12'b101010010000; // [0.66015625]
	storage[485] =  12'b101010010000; // [0.66015625]
	storage[486] =  12'b101001110000; // [0.65234375]
	storage[487] =  12'b100101010000; // [0.58203125]
	storage[488] =  12'b011100110000; // [0.44921875]
	storage[489] =  12'b010111000000; // [0.359375]
	storage[490] =  12'b010011110000; // [0.30859375]
	storage[491] =  12'b010010010000; // [0.28515625]
	storage[492] =  12'b010010100000; // [0.2890625]
	storage[493] =  12'b010100010000; // [0.31640625]
	storage[494] =  12'b010111100000; // [0.3671875]
	storage[495] =  12'b011100100000; // [0.4453125]
	storage[496] =  12'b100011100000; // [0.5546875]
	storage[497] =  12'b100111010000; // [0.61328125]
	storage[498] =  12'b101000100000; // [0.6328125]
	storage[499] =  12'b101000100000; // [0.6328125]
	storage[500] =  12'b101000010000; // [0.62890625]
	storage[501] =  12'b101000000000; // [0.625]
	storage[502] =  12'b100111110000; // [0.62109375]
	storage[503] =  12'b100111010000; // [0.61328125]
	storage[504] =  12'b100110000000; // [0.59375]
	storage[505] =  12'b100110100000; // [0.6015625]
	storage[506] =  12'b100111010000; // [0.61328125]
	storage[507] =  12'b101000000000; // [0.625]
	storage[508] =  12'b101000010000; // [0.62890625]
	storage[509] =  12'b101000110000; // [0.63671875]
	storage[510] =  12'b101001010000; // [0.64453125]
	storage[511] =  12'b101001100000; // [0.6484375]
	storage[512] =  12'b101010000000; // [0.65625]
	storage[513] =  12'b101010000000; // [0.65625]
	storage[514] =  12'b101010000000; // [0.65625]
	storage[515] =  12'b100111010000; // [0.61328125]
	storage[516] =  12'b100000110000; // [0.51171875]
	storage[517] =  12'b011001100000; // [0.3984375]
	storage[518] =  12'b010100010000; // [0.31640625]
	storage[519] =  12'b010010010000; // [0.28515625]
	storage[520] =  12'b010110000000; // [0.34375]
	storage[521] =  12'b011101010000; // [0.45703125]
	storage[522] =  12'b100010000000; // [0.53125]
	storage[523] =  12'b100100100000; // [0.5703125]
	storage[524] =  12'b100111000000; // [0.609375]
	storage[525] =  12'b101000000000; // [0.625]
	storage[526] =  12'b101000000000; // [0.625]
	storage[527] =  12'b101000000000; // [0.625]
	storage[528] =  12'b100111110000; // [0.62109375]
	storage[529] =  12'b100111100000; // [0.6171875]
	storage[530] =  12'b100111010000; // [0.61328125]
	storage[531] =  12'b100111000000; // [0.609375]
	storage[532] =  12'b100101110000; // [0.58984375]
	storage[533] =  12'b100110100000; // [0.6015625]
	storage[534] =  12'b100111000000; // [0.609375]
	storage[535] =  12'b100111110000; // [0.62109375]
	storage[536] =  12'b101000000000; // [0.625]
	storage[537] =  12'b101000110000; // [0.63671875]
	storage[538] =  12'b101001000000; // [0.640625]
	storage[539] =  12'b101001100000; // [0.6484375]
	storage[540] =  12'b101001110000; // [0.65234375]
	storage[541] =  12'b101010000000; // [0.65625]
	storage[542] =  12'b101001110000; // [0.65234375]
	storage[543] =  12'b101000100000; // [0.6328125]
	storage[544] =  12'b100101100000; // [0.5859375]
	storage[545] =  12'b011111100000; // [0.4921875]
	storage[546] =  12'b010111010000; // [0.36328125]
	storage[547] =  12'b010101010000; // [0.33203125]
	storage[548] =  12'b011011100000; // [0.4296875]
	storage[549] =  12'b100011000000; // [0.546875]
	storage[550] =  12'b100110100000; // [0.6015625]
	storage[551] =  12'b100111100000; // [0.6171875]
	storage[552] =  12'b101000000000; // [0.625]
	storage[553] =  12'b101000000000; // [0.625]
	storage[554] =  12'b101000000000; // [0.625]
	storage[555] =  12'b100111110000; // [0.62109375]
	storage[556] =  12'b100111100000; // [0.6171875]
	storage[557] =  12'b100111010000; // [0.61328125]
	storage[558] =  12'b100111000000; // [0.609375]
	storage[559] =  12'b100110100000; // [0.6015625]
	storage[560] =  12'b100101110000; // [0.58984375]
	storage[561] =  12'b100110100000; // [0.6015625]
	storage[562] =  12'b100111000000; // [0.609375]
	storage[563] =  12'b100111100000; // [0.6171875]
	storage[564] =  12'b101000000000; // [0.625]
	storage[565] =  12'b101000010000; // [0.62890625]
	storage[566] =  12'b101000110000; // [0.63671875]
	storage[567] =  12'b101001000000; // [0.640625]
	storage[568] =  12'b101001010000; // [0.64453125]
	storage[569] =  12'b101001100000; // [0.6484375]
	storage[570] =  12'b101001100000; // [0.6484375]
	storage[571] =  12'b101000000000; // [0.625]
	storage[572] =  12'b100100100000; // [0.5703125]
	storage[573] =  12'b011100000000; // [0.4375]
	storage[574] =  12'b010101100000; // [0.3359375]
	storage[575] =  12'b010111110000; // [0.37109375]
	storage[576] =  12'b011111110000; // [0.49609375]
	storage[577] =  12'b100110000000; // [0.59375]
	storage[578] =  12'b100111110000; // [0.62109375]
	storage[579] =  12'b101000010000; // [0.62890625]
	storage[580] =  12'b101000010000; // [0.62890625]
	storage[581] =  12'b101000010000; // [0.62890625]
	storage[582] =  12'b101000000000; // [0.625]
	storage[583] =  12'b100111110000; // [0.62109375]
	storage[584] =  12'b100111010000; // [0.61328125]
	storage[585] =  12'b100111000000; // [0.609375]
	storage[586] =  12'b100110110000; // [0.60546875]
	storage[587] =  12'b100110000000; // [0.59375]
	storage[588] =  12'b100101100000; // [0.5859375]
	storage[589] =  12'b100110000000; // [0.59375]
	storage[590] =  12'b100110100000; // [0.6015625]
	storage[591] =  12'b100111000000; // [0.609375]
	storage[592] =  12'b100111100000; // [0.6171875]
	storage[593] =  12'b100111110000; // [0.62109375]
	storage[594] =  12'b101000010000; // [0.62890625]
	storage[595] =  12'b101000110000; // [0.63671875]
	storage[596] =  12'b101001000000; // [0.640625]
	storage[597] =  12'b101001000000; // [0.640625]
	storage[598] =  12'b101000110000; // [0.63671875]
	storage[599] =  12'b100110110000; // [0.60546875]
	storage[600] =  12'b100001010000; // [0.51953125]
	storage[601] =  12'b011000000000; // [0.375]
	storage[602] =  12'b010101100000; // [0.3359375]
	storage[603] =  12'b011011000000; // [0.421875]
	storage[604] =  12'b100011000000; // [0.546875]
	storage[605] =  12'b100111000000; // [0.609375]
	storage[606] =  12'b101000010000; // [0.62890625]
	storage[607] =  12'b101000100000; // [0.6328125]
	storage[608] =  12'b101000100000; // [0.6328125]
	storage[609] =  12'b101000000000; // [0.625]
	storage[610] =  12'b100111100000; // [0.6171875]
	storage[611] =  12'b100111010000; // [0.61328125]
	storage[612] =  12'b100111000000; // [0.609375]
	storage[613] =  12'b100110110000; // [0.60546875]
	storage[614] =  12'b100110010000; // [0.59765625]
	storage[615] =  12'b100101110000; // [0.58984375]
	storage[616] =  12'b100101100000; // [0.5859375]
	storage[617] =  12'b100110000000; // [0.59375]
	storage[618] =  12'b100110100000; // [0.6015625]
	storage[619] =  12'b100111000000; // [0.609375]
	storage[620] =  12'b100111010000; // [0.61328125]
	storage[621] =  12'b100111100000; // [0.6171875]
	storage[622] =  12'b101000000000; // [0.625]
	storage[623] =  12'b101000010000; // [0.62890625]
	storage[624] =  12'b101000100000; // [0.6328125]
	storage[625] =  12'b101000110000; // [0.63671875]
	storage[626] =  12'b101000000000; // [0.625]
	storage[627] =  12'b100101010000; // [0.58203125]
	storage[628] =  12'b011101110000; // [0.46484375]
	storage[629] =  12'b010101100000; // [0.3359375]
	storage[630] =  12'b010110000000; // [0.34375]
	storage[631] =  12'b011101110000; // [0.46484375]
	storage[632] =  12'b100101010000; // [0.58203125]
	storage[633] =  12'b100111100000; // [0.6171875]
	storage[634] =  12'b101000010000; // [0.62890625]
	storage[635] =  12'b101000100000; // [0.6328125]
	storage[636] =  12'b101000010000; // [0.62890625]
	storage[637] =  12'b100111110000; // [0.62109375]
	storage[638] =  12'b100111100000; // [0.6171875]
	storage[639] =  12'b100111010000; // [0.61328125]
	storage[640] =  12'b100110110000; // [0.60546875]
	storage[641] =  12'b100110100000; // [0.6015625]
	storage[642] =  12'b100110000000; // [0.59375]
	storage[643] =  12'b100101100000; // [0.5859375]
	storage[644] =  12'b100101010000; // [0.58203125]
	storage[645] =  12'b100101110000; // [0.58984375]
	storage[646] =  12'b100110010000; // [0.59765625]
	storage[647] =  12'b100110100000; // [0.6015625]
	storage[648] =  12'b100111000000; // [0.609375]
	storage[649] =  12'b100111010000; // [0.61328125]
	storage[650] =  12'b100111100000; // [0.6171875]
	storage[651] =  12'b100111110000; // [0.62109375]
	storage[652] =  12'b101000000000; // [0.625]
	storage[653] =  12'b101000000000; // [0.625]
	storage[654] =  12'b100110110000; // [0.60546875]
	storage[655] =  12'b100010110000; // [0.54296875]
	storage[656] =  12'b011001100000; // [0.3984375]
	storage[657] =  12'b010100100000; // [0.3203125]
	storage[658] =  12'b010111100000; // [0.3671875]
	storage[659] =  12'b100000100000; // [0.5078125]
	storage[660] =  12'b100110010000; // [0.59765625]
	storage[661] =  12'b100111110000; // [0.62109375]
	storage[662] =  12'b101000000000; // [0.625]
	storage[663] =  12'b101000010000; // [0.62890625]
	storage[664] =  12'b101000000000; // [0.625]
	storage[665] =  12'b100111110000; // [0.62109375]
	storage[666] =  12'b100111100000; // [0.6171875]
	storage[667] =  12'b100111000000; // [0.609375]
	storage[668] =  12'b100110110000; // [0.60546875]
	storage[669] =  12'b100110010000; // [0.59765625]
	storage[670] =  12'b100101110000; // [0.58984375]
	storage[671] =  12'b100101010000; // [0.58203125]
	storage[672] =  12'b100101000000; // [0.578125]
	storage[673] =  12'b100101000000; // [0.578125]
	storage[674] =  12'b100101100000; // [0.5859375]
	storage[675] =  12'b100110000000; // [0.59375]
	storage[676] =  12'b100110100000; // [0.6015625]
	storage[677] =  12'b100110110000; // [0.60546875]
	storage[678] =  12'b100111000000; // [0.609375]
	storage[679] =  12'b100111010000; // [0.61328125]
	storage[680] =  12'b100111010000; // [0.61328125]
	storage[681] =  12'b100111010000; // [0.61328125]
	storage[682] =  12'b100101100000; // [0.5859375]
	storage[683] =  12'b011111110000; // [0.49609375]
	storage[684] =  12'b010110010000; // [0.34765625]
	storage[685] =  12'b010100000000; // [0.3125]
	storage[686] =  12'b011010000000; // [0.40625]
	storage[687] =  12'b100010110000; // [0.54296875]
	storage[688] =  12'b100111000000; // [0.609375]
	storage[689] =  12'b100111110000; // [0.62109375]
	storage[690] =  12'b101000000000; // [0.625]
	storage[691] =  12'b100111110000; // [0.62109375]
	storage[692] =  12'b100111100000; // [0.6171875]
	storage[693] =  12'b100111010000; // [0.61328125]
	storage[694] =  12'b100111000000; // [0.609375]
	storage[695] =  12'b100110110000; // [0.60546875]
	storage[696] =  12'b100110010000; // [0.59765625]
	storage[697] =  12'b100101110000; // [0.58984375]
	storage[698] =  12'b100101100000; // [0.5859375]
	storage[699] =  12'b100100110000; // [0.57421875]
	storage[700] =  12'b100100010000; // [0.56640625]
	storage[701] =  12'b100100100000; // [0.5703125]
	storage[702] =  12'b100101010000; // [0.58203125]
	storage[703] =  12'b100101110000; // [0.58984375]
	storage[704] =  12'b100110010000; // [0.59765625]
	storage[705] =  12'b100110100000; // [0.6015625]
	storage[706] =  12'b100110110000; // [0.60546875]
	storage[707] =  12'b100111000000; // [0.609375]
	storage[708] =  12'b100111000000; // [0.609375]
	storage[709] =  12'b100110110000; // [0.60546875]
	storage[710] =  12'b100100010000; // [0.56640625]
	storage[711] =  12'b011100110000; // [0.44921875]
	storage[712] =  12'b010100010000; // [0.31640625]
	storage[713] =  12'b010100100000; // [0.3203125]
	storage[714] =  12'b011100100000; // [0.4453125]
	storage[715] =  12'b100100110000; // [0.57421875]
	storage[716] =  12'b100110110000; // [0.60546875]
	storage[717] =  12'b100111010000; // [0.61328125]
	storage[718] =  12'b100111100000; // [0.6171875]
	storage[719] =  12'b100111000000; // [0.609375]
	storage[720] =  12'b100111000000; // [0.609375]
	storage[721] =  12'b100110110000; // [0.60546875]
	storage[722] =  12'b100110100000; // [0.6015625]
	storage[723] =  12'b100110010000; // [0.59765625]
	storage[724] =  12'b100110000000; // [0.59375]
	storage[725] =  12'b100101110000; // [0.58984375]
	storage[726] =  12'b100101000000; // [0.578125]
	storage[727] =  12'b100100100000; // [0.5703125]
	storage[728] =  12'b100011110000; // [0.55859375]
	storage[729] =  12'b100100010000; // [0.56640625]
	storage[730] =  12'b100101000000; // [0.578125]
	storage[731] =  12'b100101010000; // [0.58203125]
	storage[732] =  12'b100101110000; // [0.58984375]
	storage[733] =  12'b100110000000; // [0.59375]
	storage[734] =  12'b100110010000; // [0.59765625]
	storage[735] =  12'b100110010000; // [0.59765625]
	storage[736] =  12'b100110100000; // [0.6015625]
	storage[737] =  12'b100101110000; // [0.58984375]
	storage[738] =  12'b100010110000; // [0.54296875]
	storage[739] =  12'b011001100000; // [0.3984375]
	storage[740] =  12'b010011110000; // [0.30859375]
	storage[741] =  12'b010110100000; // [0.3515625]
	storage[742] =  12'b100000000000; // [0.5]
	storage[743] =  12'b100101100000; // [0.5859375]
	storage[744] =  12'b100111000000; // [0.609375]
	storage[745] =  12'b100111000000; // [0.609375]
	storage[746] =  12'b100111000000; // [0.609375]
	storage[747] =  12'b100110110000; // [0.60546875]
	storage[748] =  12'b100110110000; // [0.60546875]
	storage[749] =  12'b100110100000; // [0.6015625]
	storage[750] =  12'b100110010000; // [0.59765625]
	storage[751] =  12'b100110000000; // [0.59375]
	storage[752] =  12'b100101100000; // [0.5859375]
	storage[753] =  12'b100101000000; // [0.578125]
	storage[754] =  12'b100100110000; // [0.57421875]
	storage[755] =  12'b100100000000; // [0.5625]
	storage[756] =  12'b100010110000; // [0.54296875]
	storage[757] =  12'b100011110000; // [0.55859375]
	storage[758] =  12'b100100010000; // [0.56640625]
	storage[759] =  12'b100100110000; // [0.57421875]
	storage[760] =  12'b100101010000; // [0.58203125]
	storage[761] =  12'b100101010000; // [0.58203125]
	storage[762] =  12'b100101100000; // [0.5859375]
	storage[763] =  12'b100101110000; // [0.58984375]
	storage[764] =  12'b100101110000; // [0.58984375]
	storage[765] =  12'b100101010000; // [0.58203125]
	storage[766] =  12'b100001110000; // [0.52734375]
	storage[767] =  12'b011000110000; // [0.38671875]
	storage[768] =  12'b010100110000; // [0.32421875]
	storage[769] =  12'b011010010000; // [0.41015625]
	storage[770] =  12'b100010100000; // [0.5390625]
	storage[771] =  12'b100101110000; // [0.58984375]
	storage[772] =  12'b100110010000; // [0.59765625]
	storage[773] =  12'b100110100000; // [0.6015625]
	storage[774] =  12'b100110010000; // [0.59765625]
	storage[775] =  12'b100110010000; // [0.59765625]
	storage[776] =  12'b100110000000; // [0.59375]
	storage[777] =  12'b100110000000; // [0.59375]
	storage[778] =  12'b100101100000; // [0.5859375]
	storage[779] =  12'b100101000000; // [0.578125]
	storage[780] =  12'b100100110000; // [0.57421875]
	storage[781] =  12'b100100010000; // [0.56640625]
	storage[782] =  12'b100100000000; // [0.5625]
	storage[783] =  12'b100011010000; // [0.55078125]
end
endmodule